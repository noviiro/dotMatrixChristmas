ledmatrix
R5 7 13 100
R7 10 25 100
R3 5 15 100
R1 3 22 100
R4 6 20 100
R6 8 24 100
R2 4 16 100
R8 9 26 100

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
